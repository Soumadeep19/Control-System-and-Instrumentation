V1    1  0  PWL(0S  0V   1NS   1V   1US   1V)
R1    1  2  1KOHM
C1    2  0  1UF
.TRAN   0.1UF   10MS
.PROBE
.END
